module fetch (#parameter W=16, SIZE=20)(clk, rst, Rdst_D, Rdst_E, WD, BRANCH, FLUSH, PC_ENB, POP_L_H, JUMP_SEL, instr, imm, pc, pc_1);
    
    localparam START_ADDRESS = 2**5; //initial value of pc
    localparam ISR = 32'b0; //interrupt service routine address
    localparam NOP = 16'b0;

    input clk, rst, BRANCH, FLUSH, PC_ENB;
    input [1:0] JUMP_SEL, POP_L_H;
    input [W-1:0] Rdst_D, Rdst_E, WD;

    output [5:0] opcode;
    output [2:0] src, dst;
    output [3:0] shamt;
    output [W-1:0] instr, imm;
    output [2*W-1:0] pc, pc_1;

    reg [W-1:0] memoinst[2**SIZE-1:0];

    wire [2:0] pc_select;
    wire [2*W-1:0] ret_address, pop_in; 

    initial $readmemb("memory.txt", memoinst);

    assign pc_select = BRANCH? 3'b100: {1'b0, JUMP_SEL};

    //A temp register is used to buffer the popped address on two cycles.
    //The higher word is padded with 0's while the lower word is concatenated with the higher
    //The most significant bit in POP_L_H acts as an enable while the least
    //determines which word will be written.
    assign  pop_in = (POP_L_H == 1)? {WD, 16'b0}: {ret_address[31:16], WD}
    Register #(2*W) pc_pop (clk, rst, POP_L_H[1], pop_in, ret_address);

    mux #(2*W, 3) pc_mux ({pc+1, Rdst_D, ISR, ret_address, Rdst_E}, pc_select, pc_in)

    Register #(2*W, START_ADDRESS) pc_inst(clk, rst, PC_ENB, pc_in, pc);

    assign pc_1 = pc+1;

    assign instr = (FLUSH || BRANCH)? NOP: memoinst[pc];
    assign imm = memoinst[pc];

endmodule

//pc_sel:
// 000 pc+1
// 001 call,unconditional jump(Rdst_D)
// 010 interrupt
// 011 ret
// 100 branch(Rdst_E)
