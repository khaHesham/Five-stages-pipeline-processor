module Branch ();
    
endmodule